
module v_bb_model(CLK, STALL, RST, OPCH, OPS, TEST, AB, BC, CD, ERR, REQ, ACK, BUSY, DONE, DATA);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire [3:0] _053_;
  wire [3:0] _054_;
  wire [2:0] _055_;
  wire [2:0] _056_;
  wire [2:0] _057_;
  wire [2:0] _058_;
  output AB;
  wire AB;
  output ACK;
  reg ACK;
  output BC;
  wire BC;
  output BUSY;
  wire BUSY;
  output CD;
  wire CD;
  input CLK;
  wire CLK;
  output [2:0] DATA;
  reg [2:0] DATA;
  output DONE;
  reg DONE;
  output ERR;
  wire ERR;
  input OPCH;
  wire OPCH;
  output [3:0] OPS;
  wire [3:0] OPS;
  input REQ;
  wire REQ;
  input RST;
  wire RST;
  input STALL;
  wire STALL;
  output TEST;
  wire TEST;
  wire ack_next;
  reg [3:0] cnt;
  reg [4:0] state_reg;
  reg [2:0] unacked_reqs;
  assign _057_[0] = ~unacked_reqs[0];
  assign _053_[0] = ~cnt[0];
  assign _005_ = STALL ? state_reg[4] : state_reg[0];
  assign _015_ = state_reg[3] | state_reg[2];
  assign _002_ = STALL ? state_reg[1] : _015_;
  assign _016_ = STALL & state_reg[3];
  assign _017_ = STALL | ~(OPCH);
  assign _018_ = state_reg[4] & ~(_017_);
  assign _004_ = _018_ | _016_;
  assign _019_ = ~unacked_reqs[2];
  assign _020_ = unacked_reqs[1] | unacked_reqs[0];
  assign _021_ = _019_ & ~(_020_);
  assign _022_ = ~(cnt[1] & cnt[3]);
  assign _023_ = cnt[1] & cnt[2];
  assign _024_ = _022_ & ~(_023_);
  assign _025_ = ~(_024_ | _021_);
  assign _026_ = unacked_reqs[1] | ~(unacked_reqs[0]);
  assign _027_ = _026_ | _019_;
  assign _028_ = REQ & ~(_027_);
  assign ack_next = _028_ | _025_;
  assign _006_ = ack_next ^ REQ;
  assign _029_ = STALL & state_reg[2];
  assign _030_ = STALL | OPCH;
  assign _031_ = state_reg[4] & ~(_030_);
  assign _003_ = _031_ | _029_;
  assign _001_ = STALL ? state_reg[0] : state_reg[1];
  assign _032_ = ~(cnt[1] | cnt[0]);
  assign _033_ = ~(cnt[3] | cnt[2]);
  assign TEST = _033_ & _032_;
  assign _034_ = cnt[1] & cnt[0];
  assign _035_ = ~(cnt[3] & cnt[2]);
  assign CD = _034_ & ~(_035_);
  assign _036_ = _026_ | unacked_reqs[2];
  assign _037_ = _036_ | REQ;
  assign _000_ = ack_next & ~(_037_);
  assign _038_ = cnt[0] & ~(cnt[1]);
  assign _039_ = _038_ & _033_;
  assign _040_ = cnt[0] | ~(cnt[1]);
  assign _041_ = _033_ & ~(_040_);
  assign _042_ = _041_ | _039_;
  assign _043_ = _034_ & _033_;
  assign AB = _043_ | _042_;
  assign _044_ = cnt[3] | ~(cnt[2]);
  assign _045_ = _034_ & ~(_044_);
  assign _046_ = cnt[2] | ~(cnt[3]);
  assign _047_ = _038_ & ~(_046_);
  assign _048_ = _047_ | _045_;
  assign _049_ = _032_ & ~(_035_);
  assign BC = _049_ | _048_;
  assign BUSY = ~(_021_ | DONE);
  assign _050_ = ~(state_reg[1] | state_reg[2]);
  assign _051_ = state_reg[4] | state_reg[3];
  assign _052_ = _050_ & ~(_051_);
  assign OPS[0] = state_reg[4] & ~(_052_);
  assign OPS[1] = state_reg[3] & ~(_052_);
  assign OPS[2] = state_reg[2] & ~(_052_);
  assign OPS[3] = state_reg[1] & ~(_052_);
  assign _055_[0] = ~DATA[0];
  assign _056_[1] = DATA[1] ^ DATA[0];
  assign _007_ = DATA[1] & DATA[0];
  assign _056_[2] = _007_ ^ DATA[2];
  assign _008_ = REQ & ~(ack_next);
  assign _009_ = _008_ ^ unacked_reqs[1];
  assign _058_[1] = _009_ ^ _057_[0];
  assign _010_ = _008_ ^ unacked_reqs[2];
  assign _011_ = _008_ | ~(unacked_reqs[1]);
  assign _012_ = unacked_reqs[0] & ~(_009_);
  assign _013_ = _011_ & ~(_012_);
  assign _058_[2] = _013_ ^ _010_;
  assign _054_[1] = _038_ | ~(_040_);
  assign _054_[2] = _034_ ^ cnt[2];
  assign _014_ = _034_ & cnt[2];
  assign _054_[3] = _014_ ^ cnt[3];
  always @(posedge CLK, posedge RST)
    if (RST) DATA[0] <= 1'h0;
    else if (!ack_next) DATA[0] <= _055_[0];
  always @(posedge CLK, posedge RST)
    if (RST) DATA[1] <= 1'h0;
    else if (!ack_next) DATA[1] <= _056_[1];
  always @(posedge CLK, posedge RST)
    if (RST) DATA[2] <= 1'h0;
    else if (!ack_next) DATA[2] <= _056_[2];
  always @(posedge CLK, posedge RST)
    if (RST) state_reg[0] <= 1'h1;
    else state_reg[0] <= _001_;
  always @(posedge CLK, posedge RST)
    if (RST) state_reg[1] <= 1'h0;
    else state_reg[1] <= _002_;
  always @(posedge CLK, posedge RST)
    if (RST) state_reg[2] <= 1'h0;
    else state_reg[2] <= _003_;
  always @(posedge CLK, posedge RST)
    if (RST) state_reg[3] <= 1'h0;
    else state_reg[3] <= _004_;
  always @(posedge CLK, posedge RST)
    if (RST) state_reg[4] <= 1'h0;
    else state_reg[4] <= _005_;
  always @(posedge CLK, posedge RST)
    if (RST) unacked_reqs[0] <= 1'h0;
    else if (_006_) unacked_reqs[0] <= _057_[0];
  always @(posedge CLK, posedge RST)
    if (RST) unacked_reqs[1] <= 1'h0;
    else if (_006_) unacked_reqs[1] <= _058_[1];
  always @(posedge CLK, posedge RST)
    if (RST) unacked_reqs[2] <= 1'h0;
    else if (_006_) unacked_reqs[2] <= _058_[2];
  always @(posedge CLK, posedge RST)
    if (RST) ACK <= 1'h0;
    else ACK <= ack_next;
  always @(posedge CLK, posedge RST)
    if (RST) DONE <= 1'h0;
    else DONE <= _000_;
  always @(posedge CLK, posedge RST)
    if (RST) cnt[0] <= 1'h0;
    else cnt[0] <= _053_[0];
  always @(posedge CLK, posedge RST)
    if (RST) cnt[1] <= 1'h0;
    else cnt[1] <= _054_[1];
  always @(posedge CLK, posedge RST)
    if (RST) cnt[2] <= 1'h0;
    else cnt[2] <= _054_[2];
  always @(posedge CLK, posedge RST)
    if (RST) cnt[3] <= 1'h0;
    else cnt[3] <= _054_[3];
  assign _053_[3:1] = cnt[3:1];
  assign _054_[0] = _053_[0];
  assign _055_[2:1] = DATA[2:1];
  assign _056_[0] = _055_[0];
  assign _058_[0] = _057_[0];
  assign ERR = 1'h0;
endmodule
